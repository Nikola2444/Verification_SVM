/*******************************************************************************
    +-+-+-+-+-+-+-+-+-+-+ +-+-+-+-+-+-+-+-+-+-+-+-+ +-+-+ +-+-+-+-+-+-+-+-+
    |F|u|n|c|t|i|o|n|a|l| |V|e|r|i|f|i|c|a|t|i|o|n| |o|f| |H|a|r|d|w|a|r|e|
    +-+-+-+-+-+-+-+-+-+-+ +-+-+-+-+-+-+-+-+-+-+-+-+ +-+-+ +-+-+-+-+-+-+-+-+

    FILE            svm_dskw_seq_lib.sv

    DESCRIPTION     includes all sequences

*******************************************************************************/

//`include "sequences/svm_dskw_base_seq.sv"
`include "sequences/svm_dskw_axil_base_seq.sv"
`include "sequences/svm_dskw_axis_base_seq.sv"
`include "sequences/svm_dskw_bram_base_seq.sv"
//`include "sequences/svm_dskw_simple_seq.sv"
`include "sequences/svm_dskw_axil_seq.sv"
`include "sequences/svm_dskw_axis_seq.sv"
`include "sequences/svm_dskw_bram_seq.sv"
