Nikola@WIN-95P3O34FEFS.2196:1533981733